`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/02/01 09:32:54
// Design Name: 
// Module Name: crc_pro
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module crc_pro(
	input clk_in,
	input rst_in,
	
	input head_flag,
	input gtcrc_last_en,
	input [2:0] gtx_cnt_reside,
	input gtx_850rx_vld,
	input [63:0] gtx_850rx_dat,
	output [15:0] crc_out
    );
	
	reg [15:0] crc_buf;
	wire [63:0] d;
	wire [31:0] d_head;
	wire [7:0] d1;
	wire [15:0] d2;
	wire [23:0] d3;
	wire [31:0] d4;
	wire [39:0] d5;
	wire [47:0] d6;
	wire [55:0] d7;
	wire [15:0] c;
	
	assign d = gtx_850rx_dat;
	assign d_head = gtx_850rx_dat[31:0];
	assign d1 = gtx_850rx_dat[63:56];
	assign d2 = gtx_850rx_dat[63:48];
	assign d3 = gtx_850rx_dat[63:40];
	assign d4 = gtx_850rx_dat[63:32];
	assign d5 = gtx_850rx_dat[63:24];
	assign d6 = gtx_850rx_dat[63:16];
	assign d7 = gtx_850rx_dat[63:8];
	assign c = crc_buf;
	assign crc_out = crc_buf;
	
	always @ (posedge clk_in) begin
		if(rst_in) begin
			crc_buf <= 16'h0;
		end
		else begin
			if(gtx_850rx_vld & head_flag) begin
				crc_buf[0] <= d_head[31] ^ d_head[30] ^ d_head[27] ^ d_head[26] ^ d_head[25] ^ d_head[24] ^ d_head[23] ^ d_head[22] ^ d_head[21] ^ d_head[20] ^ d_head[19] ^ d_head[18] ^ d_head[17] ^ d_head[16] ^ d_head[15] ^ d_head[13] ^ d_head[12] ^ d_head[11] ^ d_head[10] ^ d_head[9] ^ d_head[8] ^ d_head[7] ^ d_head[6] ^ d_head[5] ^ d_head[4] ^ d_head[3] ^ d_head[2] ^ d_head[1] ^ d_head[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[14] ^ c[15];
				crc_buf[1] <= d_head[31] ^ d_head[28] ^ d_head[27] ^ d_head[26] ^ d_head[25] ^ d_head[24] ^ d_head[23] ^ d_head[22] ^ d_head[21] ^ d_head[20] ^ d_head[19] ^ d_head[18] ^ d_head[17] ^ d_head[16] ^ d_head[14] ^ d_head[13] ^ d_head[12] ^ d_head[11] ^ d_head[10] ^ d_head[9] ^ d_head[8] ^ d_head[7] ^ d_head[6] ^ d_head[5] ^ d_head[4] ^ d_head[3] ^ d_head[2] ^ d_head[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[15];
				crc_buf[2] <= d_head[31] ^ d_head[30] ^ d_head[29] ^ d_head[28] ^ d_head[16] ^ d_head[14] ^ d_head[1] ^ d_head[0] ^ c[0] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
				crc_buf[3] <= d_head[31] ^ d_head[30] ^ d_head[29] ^ d_head[17] ^ d_head[15] ^ d_head[2] ^ d_head[1] ^ c[1] ^ c[13] ^ c[14] ^ c[15];
				crc_buf[4] <= d_head[31] ^ d_head[30] ^ d_head[18] ^ d_head[16] ^ d_head[3] ^ d_head[2] ^ c[0] ^ c[2] ^ c[14] ^ c[15];
				crc_buf[5] <= d_head[31] ^ d_head[19] ^ d_head[17] ^ d_head[4] ^ d_head[3] ^ c[1] ^ c[3] ^ c[15];
				crc_buf[6] <= d_head[20] ^ d_head[18] ^ d_head[5] ^ d_head[4] ^ c[2] ^ c[4];
				crc_buf[7] <= d_head[21] ^ d_head[19] ^ d_head[6] ^ d_head[5] ^ c[3] ^ c[5];
				crc_buf[8] <= d_head[22] ^ d_head[20] ^ d_head[7] ^ d_head[6] ^ c[4] ^ c[6];
				crc_buf[9] <= d_head[23] ^ d_head[21] ^ d_head[8] ^ d_head[7] ^ c[5] ^ c[7];
				crc_buf[10] <= d_head[24] ^ d_head[22] ^ d_head[9] ^ d_head[8] ^ c[6] ^ c[8];
				crc_buf[11] <= d_head[25] ^ d_head[23] ^ d_head[10] ^ d_head[9] ^ c[7] ^ c[9];
				crc_buf[12] <= d_head[26] ^ d_head[24] ^ d_head[11] ^ d_head[10] ^ c[8] ^ c[10];
				crc_buf[13] <= d_head[27] ^ d_head[25] ^ d_head[12] ^ d_head[11] ^ c[9] ^ c[11];
				crc_buf[14] <= d_head[28] ^ d_head[26] ^ d_head[13] ^ d_head[12] ^ c[10] ^ c[12];
				crc_buf[15] <= d_head[31] ^ d_head[30] ^ d_head[29] ^ d_head[26] ^ d_head[25] ^ d_head[24] ^ d_head[23] ^ d_head[22] ^ d_head[21] ^ d_head[20] ^ d_head[19] ^ d_head[18] ^ d_head[17] ^ d_head[16] ^ d_head[15] ^ d_head[14] ^ d_head[12] ^ d_head[11] ^ d_head[10] ^ d_head[9] ^ d_head[8] ^ d_head[7] ^ d_head[6] ^ d_head[5] ^ d_head[4] ^ d_head[3] ^ d_head[2] ^ d_head[1] ^ d_head[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[15];
			end
			else if(gtx_850rx_vld & gtcrc_last_en) begin
				case(gtx_cnt_reside)
					3'd1: begin
						crc_buf[0] <= d1[7] ^ d1[6] ^ d1[5] ^ d1[4] ^ d1[3] ^ d1[2] ^ d1[1] ^ d1[0] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[1] <= d1[7] ^ d1[6] ^ d1[5] ^ d1[4] ^ d1[3] ^ d1[2] ^ d1[1] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[2] <= d1[1] ^ d1[0] ^ c[8] ^ c[9];
						crc_buf[3] <= d1[2] ^ d1[1] ^ c[9] ^ c[10];
						crc_buf[4] <= d1[3] ^ d1[2] ^ c[10] ^ c[11];
						crc_buf[5] <= d1[4] ^ d1[3] ^ c[11] ^ c[12];
						crc_buf[6] <= d1[5] ^ d1[4] ^ c[12] ^ c[13];
						crc_buf[7] <= d1[6] ^ d1[5] ^ c[13] ^ c[14];
						crc_buf[8] <= d1[7] ^ d1[6] ^ c[0] ^ c[14] ^ c[15];
						crc_buf[9] <= d1[7] ^ c[1] ^ c[15];
						crc_buf[10] <= c[2];
						crc_buf[11] <= c[3];
						crc_buf[12] <= c[4];
						crc_buf[13] <= c[5];
						crc_buf[14] <= c[6];
						crc_buf[15] <= d1[7] ^ d1[6] ^ d1[5] ^ d1[4] ^ d1[3] ^ d1[2] ^ d1[1] ^ d1[0] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
					end
					3'd2: begin
						crc_buf[0] <= d2[15] ^ d2[13] ^ d2[12] ^ d2[11] ^ d2[10] ^ d2[9] ^ d2[8] ^ d2[7] ^ d2[6] ^ d2[5] ^ d2[4] ^ d2[3] ^ d2[2] ^ d2[1] ^ d2[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[15];
						crc_buf[1] <= d2[14] ^ d2[13] ^ d2[12] ^ d2[11] ^ d2[10] ^ d2[9] ^ d2[8] ^ d2[7] ^ d2[6] ^ d2[5] ^ d2[4] ^ d2[3] ^ d2[2] ^ d2[1] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14];
						crc_buf[2] <= d2[14] ^ d2[1] ^ d2[0] ^ c[0] ^ c[1] ^ c[14];
						crc_buf[3] <= d2[15] ^ d2[2] ^ d2[1] ^ c[1] ^ c[2] ^ c[15];
						crc_buf[4] <= d2[3] ^ d2[2] ^ c[2] ^ c[3];
						crc_buf[5] <= d2[4] ^ d2[3] ^ c[3] ^ c[4];
						crc_buf[6] <= d2[5] ^ d2[4] ^ c[4] ^ c[5];
						crc_buf[7] <= d2[6] ^ d2[5] ^ c[5] ^ c[6];
						crc_buf[8] <= d2[7] ^ d2[6] ^ c[6] ^ c[7];
						crc_buf[9] <= d2[8] ^ d2[7] ^ c[7] ^ c[8];
						crc_buf[10] <= d2[9] ^ d2[8] ^ c[8] ^ c[9];
						crc_buf[11] <= d2[10] ^ d2[9] ^ c[9] ^ c[10];
						crc_buf[12] <= d2[11] ^ d2[10] ^ c[10] ^ c[11];
						crc_buf[13] <= d2[12] ^ d2[11] ^ c[11] ^ c[12];
						crc_buf[14] <= d2[13] ^ d2[12] ^ c[12] ^ c[13];
						crc_buf[15] <= d2[15] ^ d2[14] ^ d2[12] ^ d2[11] ^ d2[10] ^ d2[9] ^ d2[8] ^ d2[7] ^ d2[6] ^ d2[5] ^ d2[4] ^ d2[3] ^ d2[2] ^ d2[1] ^ d2[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[14] ^ c[15];
					end
					3'd3: begin
						crc_buf[0] <= d3[23] ^ d3[22] ^ d3[21] ^ d3[20] ^ d3[19] ^ d3[18] ^ d3[17] ^ d3[16] ^ d3[15] ^ d3[13] ^ d3[12] ^ d3[11] ^ d3[10] ^ d3[9] ^ d3[8] ^ d3[7] ^ d3[6] ^ d3[5] ^ d3[4] ^ d3[3] ^ d3[2] ^ d3[1] ^ d3[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[1] <= d3[23] ^ d3[22] ^ d3[21] ^ d3[20] ^ d3[19] ^ d3[18] ^ d3[17] ^ d3[16] ^ d3[14] ^ d3[13] ^ d3[12] ^ d3[11] ^ d3[10] ^ d3[9] ^ d3[8] ^ d3[7] ^ d3[6] ^ d3[5] ^ d3[4] ^ d3[3] ^ d3[2] ^ d3[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[2] <= d3[16] ^ d3[14] ^ d3[1] ^ d3[0] ^ c[6] ^ c[8];
						crc_buf[3] <= d3[17] ^ d3[15] ^ d3[2] ^ d3[1] ^ c[7] ^ c[9];
						crc_buf[4] <= d3[18] ^ d3[16] ^ d3[3] ^ d3[2] ^ c[8] ^ c[10];
						crc_buf[5] <= d3[19] ^ d3[17] ^ d3[4] ^ d3[3] ^ c[9] ^ c[11];
						crc_buf[6] <= d3[20] ^ d3[18] ^ d3[5] ^ d3[4] ^ c[10] ^ c[12];
						crc_buf[7] <= d3[21] ^ d3[19] ^ d3[6] ^ d3[5] ^ c[11] ^ c[13];
						crc_buf[8] <= d3[22] ^ d3[20] ^ d3[7] ^ d3[6] ^ c[12] ^ c[14];
						crc_buf[9] <= d3[23] ^ d3[21] ^ d3[8] ^ d3[7] ^ c[0] ^ c[13] ^ c[15];
						crc_buf[10] <= d3[22] ^ d3[9] ^ d3[8] ^ c[0] ^ c[1] ^ c[14];
						crc_buf[11] <= d3[23] ^ d3[10] ^ d3[9] ^ c[1] ^ c[2] ^ c[15];
						crc_buf[12] <= d3[11] ^ d3[10] ^ c[2] ^ c[3];
						crc_buf[13] <= d3[12] ^ d3[11] ^ c[3] ^ c[4];
						crc_buf[14] <= d3[13] ^ d3[12] ^ c[4] ^ c[5];
						crc_buf[15] <= d3[23] ^ d3[22] ^ d3[21] ^ d3[20] ^ d3[19] ^ d3[18] ^ d3[17] ^ d3[16] ^ d3[15] ^ d3[14] ^ d3[12] ^ d3[11] ^ d3[10] ^ d3[9] ^ d3[8] ^ d3[7] ^ d3[6] ^ d3[5] ^ d3[4] ^ d3[3] ^ d3[2] ^ d3[1] ^ d3[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
					end
					3'd4: begin
						crc_buf[0] <= d4[31] ^ d4[30] ^ d4[27] ^ d4[26] ^ d4[25] ^ d4[24] ^ d4[23] ^ d4[22] ^ d4[21] ^ d4[20] ^ d4[19] ^ d4[18] ^ d4[17] ^ d4[16] ^ d4[15] ^ d4[13] ^ d4[12] ^ d4[11] ^ d4[10] ^ d4[9] ^ d4[8] ^ d4[7] ^ d4[6] ^ d4[5] ^ d4[4] ^ d4[3] ^ d4[2] ^ d4[1] ^ d4[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[14] ^ c[15];
						crc_buf[1] <= d4[31] ^ d4[28] ^ d4[27] ^ d4[26] ^ d4[25] ^ d4[24] ^ d4[23] ^ d4[22] ^ d4[21] ^ d4[20] ^ d4[19] ^ d4[18] ^ d4[17] ^ d4[16] ^ d4[14] ^ d4[13] ^ d4[12] ^ d4[11] ^ d4[10] ^ d4[9] ^ d4[8] ^ d4[7] ^ d4[6] ^ d4[5] ^ d4[4] ^ d4[3] ^ d4[2] ^ d4[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[15];
						crc_buf[2] <= d4[31] ^ d4[30] ^ d4[29] ^ d4[28] ^ d4[16] ^ d4[14] ^ d4[1] ^ d4[0] ^ c[0] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[3] <= d4[31] ^ d4[30] ^ d4[29] ^ d4[17] ^ d4[15] ^ d4[2] ^ d4[1] ^ c[1] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[4] <= d4[31] ^ d4[30] ^ d4[18] ^ d4[16] ^ d4[3] ^ d4[2] ^ c[0] ^ c[2] ^ c[14] ^ c[15];
						crc_buf[5] <= d4[31] ^ d4[19] ^ d4[17] ^ d4[4] ^ d4[3] ^ c[1] ^ c[3] ^ c[15];
						crc_buf[6] <= d4[20] ^ d4[18] ^ d4[5] ^ d4[4] ^ c[2] ^ c[4];
						crc_buf[7] <= d4[21] ^ d4[19] ^ d4[6] ^ d4[5] ^ c[3] ^ c[5];
						crc_buf[8] <= d4[22] ^ d4[20] ^ d4[7] ^ d4[6] ^ c[4] ^ c[6];
						crc_buf[9] <= d4[23] ^ d4[21] ^ d4[8] ^ d4[7] ^ c[5] ^ c[7];
						crc_buf[10] <= d4[24] ^ d4[22] ^ d4[9] ^ d4[8] ^ c[6] ^ c[8];
						crc_buf[11] <= d4[25] ^ d4[23] ^ d4[10] ^ d4[9] ^ c[7] ^ c[9];
						crc_buf[12] <= d4[26] ^ d4[24] ^ d4[11] ^ d4[10] ^ c[8] ^ c[10];
						crc_buf[13] <= d4[27] ^ d4[25] ^ d4[12] ^ d4[11] ^ c[9] ^ c[11];
						crc_buf[14] <= d4[28] ^ d4[26] ^ d4[13] ^ d4[12] ^ c[10] ^ c[12];
						crc_buf[15] <= d4[31] ^ d4[30] ^ d4[29] ^ d4[26] ^ d4[25] ^ d4[24] ^ d4[23] ^ d4[22] ^ d4[21] ^ d4[20] ^ d4[19] ^ d4[18] ^ d4[17] ^ d4[16] ^ d4[15] ^ d4[14] ^ d4[12] ^ d4[11] ^ d4[10] ^ d4[9] ^ d4[8] ^ d4[7] ^ d4[6] ^ d4[5] ^ d4[4] ^ d4[3] ^ d4[2] ^ d4[1] ^ d4[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[15];
					end
					3'd5: begin
						crc_buf[0] <= d5[39] ^ d5[38] ^ d5[37] ^ d5[36] ^ d5[35] ^ d5[34] ^ d5[33] ^ d5[32] ^ d5[31] ^ d5[30] ^ d5[27] ^ d5[26] ^ d5[25] ^ d5[24] ^ d5[23] ^ d5[22] ^ d5[21] ^ d5[20] ^ d5[19] ^ d5[18] ^ d5[17] ^ d5[16] ^ d5[15] ^ d5[13] ^ d5[12] ^ d5[11] ^ d5[10] ^ d5[9] ^ d5[8] ^ d5[7] ^ d5[6] ^ d5[5] ^ d5[4] ^ d5[3] ^ d5[2] ^ d5[1] ^ d5[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[1] <= d5[39] ^ d5[38] ^ d5[37] ^ d5[36] ^ d5[35] ^ d5[34] ^ d5[33] ^ d5[32] ^ d5[31] ^ d5[28] ^ d5[27] ^ d5[26] ^ d5[25] ^ d5[24] ^ d5[23] ^ d5[22] ^ d5[21] ^ d5[20] ^ d5[19] ^ d5[18] ^ d5[17] ^ d5[16] ^ d5[14] ^ d5[13] ^ d5[12] ^ d5[11] ^ d5[10] ^ d5[9] ^ d5[8] ^ d5[7] ^ d5[6] ^ d5[5] ^ d5[4] ^ d5[3] ^ d5[2] ^ d5[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[2] <= d5[31] ^ d5[30] ^ d5[29] ^ d5[28] ^ d5[16] ^ d5[14] ^ d5[1] ^ d5[0] ^ c[4] ^ c[5] ^ c[6] ^ c[7];
						crc_buf[3] <= d5[32] ^ d5[31] ^ d5[30] ^ d5[29] ^ d5[17] ^ d5[15] ^ d5[2] ^ d5[1] ^ c[5] ^ c[6] ^ c[7] ^ c[8];
						crc_buf[4] <= d5[33] ^ d5[32] ^ d5[31] ^ d5[30] ^ d5[18] ^ d5[16] ^ d5[3] ^ d5[2] ^ c[6] ^ c[7] ^ c[8] ^ c[9];
						crc_buf[5] <= d5[34] ^ d5[33] ^ d5[32] ^ d5[31] ^ d5[19] ^ d5[17] ^ d5[4] ^ d5[3] ^ c[7] ^ c[8] ^ c[9] ^ c[10];
						crc_buf[6] <= d5[35] ^ d5[34] ^ d5[33] ^ d5[32] ^ d5[20] ^ d5[18] ^ d5[5] ^ d5[4] ^ c[8] ^ c[9] ^ c[10] ^ c[11];
						crc_buf[7] <= d5[36] ^ d5[35] ^ d5[34] ^ d5[33] ^ d5[21] ^ d5[19] ^ d5[6] ^ d5[5] ^ c[9] ^ c[10] ^ c[11] ^ c[12];
						crc_buf[8] <= d5[37] ^ d5[36] ^ d5[35] ^ d5[34] ^ d5[22] ^ d5[20] ^ d5[7] ^ d5[6] ^ c[10] ^ c[11] ^ c[12] ^ c[13];
						crc_buf[9] <= d5[38] ^ d5[37] ^ d5[36] ^ d5[35] ^ d5[23] ^ d5[21] ^ d5[8] ^ d5[7] ^ c[11] ^ c[12] ^ c[13] ^ c[14];
						crc_buf[10] <= d5[39] ^ d5[38] ^ d5[37] ^ d5[36] ^ d5[24] ^ d5[22] ^ d5[9] ^ d5[8] ^ c[0] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[11] <= d5[39] ^ d5[38] ^ d5[37] ^ d5[25] ^ d5[23] ^ d5[10] ^ d5[9] ^ c[1] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[12] <= d5[39] ^ d5[38] ^ d5[26] ^ d5[24] ^ d5[11] ^ d5[10] ^ c[0] ^ c[2] ^ c[14] ^ c[15];
						crc_buf[13] <= d5[39] ^ d5[27] ^ d5[25] ^ d5[12] ^ d5[11] ^ c[1] ^ c[3] ^ c[15];
						crc_buf[14] <= d5[28] ^ d5[26] ^ d5[13] ^ d5[12] ^ c[2] ^ c[4];
						crc_buf[15] <= d5[39] ^ d5[38] ^ d5[37] ^ d5[36] ^ d5[35] ^ d5[34] ^ d5[33] ^ d5[32] ^ d5[31] ^ d5[30] ^ d5[29] ^ d5[26] ^ d5[25] ^ d5[24] ^ d5[23] ^ d5[22] ^ d5[21] ^ d5[20] ^ d5[19] ^ d5[18] ^ d5[17] ^ d5[16] ^ d5[15] ^ d5[14] ^ d5[12] ^ d5[11] ^ d5[10] ^ d5[9] ^ d5[8] ^ d5[7] ^ d5[6] ^ d5[5] ^ d5[4] ^ d5[3] ^ d5[2] ^ d5[1] ^ d5[0] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
					end
					3'd6: begin
						crc_buf[0] <= d6[47] ^ d6[46] ^ d6[45] ^ d6[43] ^ d6[41] ^ d6[40] ^ d6[39] ^ d6[38] ^ d6[37] ^ d6[36] ^ d6[35] ^ d6[34] ^ d6[33] ^ d6[32] ^ d6[31] ^ d6[30] ^ d6[27] ^ d6[26] ^ d6[25] ^ d6[24] ^ d6[23] ^ d6[22] ^ d6[21] ^ d6[20] ^ d6[19] ^ d6[18] ^ d6[17] ^ d6[16] ^ d6[15] ^ d6[13] ^ d6[12] ^ d6[11] ^ d6[10] ^ d6[9] ^ d6[8] ^ d6[7] ^ d6[6] ^ d6[5] ^ d6[4] ^ d6[3] ^ d6[2] ^ d6[1] ^ d6[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[1] <= d6[47] ^ d6[46] ^ d6[44] ^ d6[42] ^ d6[41] ^ d6[40] ^ d6[39] ^ d6[38] ^ d6[37] ^ d6[36] ^ d6[35] ^ d6[34] ^ d6[33] ^ d6[32] ^ d6[31] ^ d6[28] ^ d6[27] ^ d6[26] ^ d6[25] ^ d6[24] ^ d6[23] ^ d6[22] ^ d6[21] ^ d6[20] ^ d6[19] ^ d6[18] ^ d6[17] ^ d6[16] ^ d6[14] ^ d6[13] ^ d6[12] ^ d6[11] ^ d6[10] ^ d6[9] ^ d6[8] ^ d6[7] ^ d6[6] ^ d6[5] ^ d6[4] ^ d6[3] ^ d6[2] ^ d6[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[14] ^ c[15];
						crc_buf[2] <= d6[46] ^ d6[42] ^ d6[31] ^ d6[30] ^ d6[29] ^ d6[28] ^ d6[16] ^ d6[14] ^ d6[1] ^ d6[0] ^ c[10] ^ c[14];
						crc_buf[3] <= d6[47] ^ d6[43] ^ d6[32] ^ d6[31] ^ d6[30] ^ d6[29] ^ d6[17] ^ d6[15] ^ d6[2] ^ d6[1] ^ c[0] ^ c[11] ^ c[15];
						crc_buf[4] <= d6[44] ^ d6[33] ^ d6[32] ^ d6[31] ^ d6[30] ^ d6[18] ^ d6[16] ^ d6[3] ^ d6[2] ^ c[0] ^ c[1] ^ c[12];
						crc_buf[5] <= d6[45] ^ d6[34] ^ d6[33] ^ d6[32] ^ d6[31] ^ d6[19] ^ d6[17] ^ d6[4] ^ d6[3] ^ c[0] ^ c[1] ^ c[2] ^ c[13];
						crc_buf[6] <= d6[46] ^ d6[35] ^ d6[34] ^ d6[33] ^ d6[32] ^ d6[20] ^ d6[18] ^ d6[5] ^ d6[4] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[14];
						crc_buf[7] <= d6[47] ^ d6[36] ^ d6[35] ^ d6[34] ^ d6[33] ^ d6[21] ^ d6[19] ^ d6[6] ^ d6[5] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[15];
						crc_buf[8] <= d6[37] ^ d6[36] ^ d6[35] ^ d6[34] ^ d6[22] ^ d6[20] ^ d6[7] ^ d6[6] ^ c[2] ^ c[3] ^ c[4] ^ c[5];
						crc_buf[9] <= d6[38] ^ d6[37] ^ d6[36] ^ d6[35] ^ d6[23] ^ d6[21] ^ d6[8] ^ d6[7] ^ c[3] ^ c[4] ^ c[5] ^ c[6];
						crc_buf[10] <= d6[39] ^ d6[38] ^ d6[37] ^ d6[36] ^ d6[24] ^ d6[22] ^ d6[9] ^ d6[8] ^ c[4] ^ c[5] ^ c[6] ^ c[7];
						crc_buf[11] <= d6[40] ^ d6[39] ^ d6[38] ^ d6[37] ^ d6[25] ^ d6[23] ^ d6[10] ^ d6[9] ^ c[5] ^ c[6] ^ c[7] ^ c[8];
						crc_buf[12] <= d6[41] ^ d6[40] ^ d6[39] ^ d6[38] ^ d6[26] ^ d6[24] ^ d6[11] ^ d6[10] ^ c[6] ^ c[7] ^ c[8] ^ c[9];
						crc_buf[13] <= d6[42] ^ d6[41] ^ d6[40] ^ d6[39] ^ d6[27] ^ d6[25] ^ d6[12] ^ d6[11] ^ c[7] ^ c[8] ^ c[9] ^ c[10];
						crc_buf[14] <= d6[43] ^ d6[42] ^ d6[41] ^ d6[40] ^ d6[28] ^ d6[26] ^ d6[13] ^ d6[12] ^ c[8] ^ c[9] ^ c[10] ^ c[11];
						crc_buf[15] <= d6[47] ^ d6[46] ^ d6[45] ^ d6[44] ^ d6[42] ^ d6[40] ^ d6[39] ^ d6[38] ^ d6[37] ^ d6[36] ^ d6[35] ^ d6[34] ^ d6[33] ^ d6[32] ^ d6[31] ^ d6[30] ^ d6[29] ^ d6[26] ^ d6[25] ^ d6[24] ^ d6[23] ^ d6[22] ^ d6[21] ^ d6[20] ^ d6[19] ^ d6[18] ^ d6[17] ^ d6[16] ^ d6[15] ^ d6[14] ^ d6[12] ^ d6[11] ^ d6[10] ^ d6[9] ^ d6[8] ^ d6[7] ^ d6[6] ^ d6[5] ^ d6[4] ^ d6[3] ^ d6[2] ^ d6[1] ^ d6[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
					end
					3'd7: begin
						crc_buf[0] <= d7[55] ^ d7[54] ^ d7[53] ^ d7[52] ^ d7[51] ^ d7[50] ^ d7[49] ^ d7[48] ^ d7[47] ^ d7[46] ^ d7[45] ^ d7[43] ^ d7[41] ^ d7[40] ^ d7[39] ^ d7[38] ^ d7[37] ^ d7[36] ^ d7[35] ^ d7[34] ^ d7[33] ^ d7[32] ^ d7[31] ^ d7[30] ^ d7[27] ^ d7[26] ^ d7[25] ^ d7[24] ^ d7[23] ^ d7[22] ^ d7[21] ^ d7[20] ^ d7[19] ^ d7[18] ^ d7[17] ^ d7[16] ^ d7[15] ^ d7[13] ^ d7[12] ^ d7[11] ^ d7[10] ^ d7[9] ^ d7[8] ^ d7[7] ^ d7[6] ^ d7[5] ^ d7[4] ^ d7[3] ^ d7[2] ^ d7[1] ^ d7[0] ^ c[0] ^ c[1] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[1] <= d7[55] ^ d7[54] ^ d7[53] ^ d7[52] ^ d7[51] ^ d7[50] ^ d7[49] ^ d7[48] ^ d7[47] ^ d7[46] ^ d7[44] ^ d7[42] ^ d7[41] ^ d7[40] ^ d7[39] ^ d7[38] ^ d7[37] ^ d7[36] ^ d7[35] ^ d7[34] ^ d7[33] ^ d7[32] ^ d7[31] ^ d7[28] ^ d7[27] ^ d7[26] ^ d7[25] ^ d7[24] ^ d7[23] ^ d7[22] ^ d7[21] ^ d7[20] ^ d7[19] ^ d7[18] ^ d7[17] ^ d7[16] ^ d7[14] ^ d7[13] ^ d7[12] ^ d7[11] ^ d7[10] ^ d7[9] ^ d7[8] ^ d7[7] ^ d7[6] ^ d7[5] ^ d7[4] ^ d7[3] ^ d7[2] ^ d7[1] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
						crc_buf[2] <= d7[46] ^ d7[42] ^ d7[31] ^ d7[30] ^ d7[29] ^ d7[28] ^ d7[16] ^ d7[14] ^ d7[1] ^ d7[0] ^ c[2] ^ c[6];
						crc_buf[3] <= d7[47] ^ d7[43] ^ d7[32] ^ d7[31] ^ d7[30] ^ d7[29] ^ d7[17] ^ d7[15] ^ d7[2] ^ d7[1] ^ c[3] ^ c[7];
						crc_buf[4] <= d7[48] ^ d7[44] ^ d7[33] ^ d7[32] ^ d7[31] ^ d7[30] ^ d7[18] ^ d7[16] ^ d7[3] ^ d7[2] ^ c[4] ^ c[8];
						crc_buf[5] <= d7[49] ^ d7[45] ^ d7[34] ^ d7[33] ^ d7[32] ^ d7[31] ^ d7[19] ^ d7[17] ^ d7[4] ^ d7[3] ^ c[5] ^ c[9];
						crc_buf[6] <= d7[50] ^ d7[46] ^ d7[35] ^ d7[34] ^ d7[33] ^ d7[32] ^ d7[20] ^ d7[18] ^ d7[5] ^ d7[4] ^ c[6] ^ c[10];
						crc_buf[7] <= d7[51] ^ d7[47] ^ d7[36] ^ d7[35] ^ d7[34] ^ d7[33] ^ d7[21] ^ d7[19] ^ d7[6] ^ d7[5] ^ c[7] ^ c[11];
						crc_buf[8] <= d7[52] ^ d7[48] ^ d7[37] ^ d7[36] ^ d7[35] ^ d7[34] ^ d7[22] ^ d7[20] ^ d7[7] ^ d7[6] ^ c[8] ^ c[12];
						crc_buf[9] <= d7[53] ^ d7[49] ^ d7[38] ^ d7[37] ^ d7[36] ^ d7[35] ^ d7[23] ^ d7[21] ^ d7[8] ^ d7[7] ^ c[9] ^ c[13];
						crc_buf[10] <= d7[54] ^ d7[50] ^ d7[39] ^ d7[38] ^ d7[37] ^ d7[36] ^ d7[24] ^ d7[22] ^ d7[9] ^ d7[8] ^ c[10] ^ c[14];
						crc_buf[11] <= d7[55] ^ d7[51] ^ d7[40] ^ d7[39] ^ d7[38] ^ d7[37] ^ d7[25] ^ d7[23] ^ d7[10] ^ d7[9] ^ c[0] ^ c[11] ^ c[15];
						crc_buf[12] <= d7[52] ^ d7[41] ^ d7[40] ^ d7[39] ^ d7[38] ^ d7[26] ^ d7[24] ^ d7[11] ^ d7[10] ^ c[0] ^ c[1] ^ c[12];
						crc_buf[13] <= d7[53] ^ d7[42] ^ d7[41] ^ d7[40] ^ d7[39] ^ d7[27] ^ d7[25] ^ d7[12] ^ d7[11] ^ c[0] ^ c[1] ^ c[2] ^ c[13];
						crc_buf[14] <= d7[54] ^ d7[43] ^ d7[42] ^ d7[41] ^ d7[40] ^ d7[28] ^ d7[26] ^ d7[13] ^ d7[12] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[14];
						crc_buf[15] <= d7[54] ^ d7[53] ^ d7[52] ^ d7[51] ^ d7[50] ^ d7[49] ^ d7[48] ^ d7[47] ^ d7[46] ^ d7[45] ^ d7[44] ^ d7[42] ^ d7[40] ^ d7[39] ^ d7[38] ^ d7[37] ^ d7[36] ^ d7[35] ^ d7[34] ^ d7[33] ^ d7[32] ^ d7[31] ^ d7[30] ^ d7[29] ^ d7[26] ^ d7[25] ^ d7[24] ^ d7[23] ^ d7[22] ^ d7[21] ^ d7[20] ^ d7[19] ^ d7[18] ^ d7[17] ^ d7[16] ^ d7[15] ^ d7[14] ^ d7[12] ^ d7[11] ^ d7[10] ^ d7[9] ^ d7[8] ^ d7[7] ^ d7[6] ^ d7[5] ^ d7[4] ^ d7[3] ^ d7[2] ^ d7[1] ^ d7[0] ^ c[0] ^ c[2] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14];
					end
				endcase
			end
			else if(gtx_850rx_vld) begin
				crc_buf[0] <= d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[13] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
				crc_buf[1] <= d[63] ^ d[62] ^ d[61] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[31] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[13] ^ c[14] ^ c[15];
				crc_buf[2] <= d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[46] ^ d[42] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[16] ^ d[14] ^ d[1] ^ d[0] ^ c[8] ^ c[9] ^ c[12] ^ c[13];
				crc_buf[3] <= d[62] ^ d[61] ^ d[58] ^ d[57] ^ d[47] ^ d[43] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[17] ^ d[15] ^ d[2] ^ d[1] ^ c[9] ^ c[10] ^ c[13] ^ c[14];
				crc_buf[4] <= d[63] ^ d[62] ^ d[59] ^ d[58] ^ d[48] ^ d[44] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[18] ^ d[16] ^ d[3] ^ d[2] ^ c[0] ^ c[10] ^ c[11] ^ c[14] ^ c[15];
				crc_buf[5] <= d[63] ^ d[60] ^ d[59] ^ d[49] ^ d[45] ^ d[34] ^ d[33] ^ d[32] ^ d[31] ^ d[19] ^ d[17] ^ d[4] ^ d[3] ^ c[1] ^ c[11] ^ c[12] ^ c[15];
				crc_buf[6] <= d[61] ^ d[60] ^ d[50] ^ d[46] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[20] ^ d[18] ^ d[5] ^ d[4] ^ c[2] ^ c[12] ^ c[13];
				crc_buf[7] <= d[62] ^ d[61] ^ d[51] ^ d[47] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[21] ^ d[19] ^ d[6] ^ d[5] ^ c[3] ^ c[13] ^ c[14];
				crc_buf[8] <= d[63] ^ d[62] ^ d[52] ^ d[48] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[22] ^ d[20] ^ d[7] ^ d[6] ^ c[0] ^ c[4] ^ c[14] ^ c[15];
				crc_buf[9] <= d[63] ^ d[53] ^ d[49] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[23] ^ d[21] ^ d[8] ^ d[7] ^ c[1] ^ c[5] ^ c[15];
				crc_buf[10] <= d[54] ^ d[50] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[24] ^ d[22] ^ d[9] ^ d[8] ^ c[2] ^ c[6];
				crc_buf[11] <= d[55] ^ d[51] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[25] ^ d[23] ^ d[10] ^ d[9] ^ c[3] ^ c[7];
				crc_buf[12] <= d[56] ^ d[52] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[26] ^ d[24] ^ d[11] ^ d[10] ^ c[4] ^ c[8];
				crc_buf[13] <= d[57] ^ d[53] ^ d[42] ^ d[41] ^ d[40] ^ d[39] ^ d[27] ^ d[25] ^ d[12] ^ d[11] ^ c[5] ^ c[9];
				crc_buf[14] <= d[58] ^ d[54] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[28] ^ d[26] ^ d[13] ^ d[12] ^ c[6] ^ c[10];
				crc_buf[15] <= d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15];
			end
			else begin
				crc_buf <= crc_buf;
			end
		end
	end
	
endmodule
